// ********************************************************************
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// ********************************************************************
// File name    : led.v
// Module name  : led
// Author       : STEP
// Description  : control LED
// Web          : www.stepfpga.com
// 
// --------------------------------------------------------------------
// Code Revision History : 
// --------------------------------------------------------------------
// Version: |Mod. Date:   |Changes Made:
// V1.0     |2017/03/02   |Initial ver
// --------------------------------------------------------------------
// Module Function:���ð����Ϳ��ص�״̬������LED�Ƶ�����
 
module led (key,sw,led);
 
	input [3:0] key;						//���������ź�
	input [3:0] sw;							//���������ź�
	output [7:0] led;						//����źŵ�LED
 
	assign led = {key,sw};                  //assign������ֵ����������ƴ�ӷ�����ʾ��key��swƴ�����һ���µ�8λ����ֵ��led
 
endmodule